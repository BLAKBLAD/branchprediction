`timescale 1ns / 1ps

module module_gshare(

    );
endmodule
